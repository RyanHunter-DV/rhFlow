// standard sv file 
