class rh_axi4_drvBase#(type REQ=rh_axi4_trans,RSP=REQ) extends uvm_driver#(REQ,RSP);
	<extra>
	`uvm_component_utils_begin(rh_axi4_drvBase)
	`uvm_component_utils_end
